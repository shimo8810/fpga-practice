module vga(
    input logic pixclk
    );
    // �g�b�v�Ƃ���
endmodule
