`ifndef LIB_VGA_SVH
`define LIB_VGA_SVH
package libvga;


endpackage
`endif